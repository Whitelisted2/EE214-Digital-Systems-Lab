	else
	   bin_out(0) <= '0';
		bin_out(1) <= '0';
	end if;
	end process c1;
end behavioral;